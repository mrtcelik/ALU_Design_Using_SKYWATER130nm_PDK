** sch_path: /home/halil/Desktop/design/xschem/8bit_multiplier.sch
**.subckt 8bit_multiplier VDD VSS A0 A1 A2 A3 B1 mult_out0 B0 mult_out1 B2 B3 mult_out2 mult_out3
*+ mult_out4 mult_out5 mult_out6 mult_out7
*.iopin VDD
*.iopin VSS
*.ipin A0
*.ipin A1
*.ipin A2
*.ipin A3
*.ipin B1
*.opin mult_out0
*.ipin B0
*.opin mult_out1
*.ipin B2
*.ipin B3
*.opin mult_out2
*.opin mult_out3
*.opin mult_out4
*.opin mult_out5
*.opin mult_out6
*.opin mult_out7
x1 VDD VSS net9 net10 net11 mult_out1 net7 net1 net8 VSS net6 net3 net4 net5 net2 4bit_adder
x2 VSS VDD A0 mult_out0 B0 and2
x3 VSS VDD A1 net1 B0 and2
x4 VSS VDD A2 net2 B0 and2
x5 VSS VDD A3 net3 B0 and2
x6 VSS VDD A0 net7 B1 and2
x7 VSS VDD A1 net4 B1 and2
x8 VSS VDD A2 net5 B1 and2
x9 VSS VDD A3 net6 B1 and2
x10 VDD VSS net18 net17 net16 mult_out2 net15 net11 net19 net8 net12 net9 net14 net13 net10
+ 4bit_adder
x11 VSS VDD A0 net15 B2 and2
x12 VSS VDD A1 net14 B2 and2
x13 VSS VDD A2 net13 B2 and2
x14 VSS VDD A3 net12 B2 and2
x15 VDD VSS mult_out6 mult_out5 mult_out4 mult_out3 net23 net16 mult_out7 net19 net20 net18 net22
+ net21 net17 4bit_adder
x16 VSS VDD A0 net23 B3 and2
x17 VSS VDD A1 net22 B3 and2
x18 VSS VDD A2 net21 B3 and2
x19 VSS VDD A3 net20 B3 and2
**.ends

* expanding   symbol:  adder/4bit_adder.sym # of pins=15
** sym_path: /home/halil/Desktop/design/xschem/adder/4bit_adder.sym
** sch_path: /home/halil/Desktop/design/xschem/adder/4bit_adder.sch
.subckt 4bit_adder  VDD VSS adder_out3 adder_out2 adder_out1 adder_out0 A0 B0 Cout B3 A3 B2 A1 A2 B1
*.iopin VDD
*.iopin VSS
*.ipin B0
*.ipin A1
*.ipin B1
*.opin adder_out0
*.ipin A2
*.ipin B2
*.opin adder_out1
*.opin adder_out2
*.ipin A3
*.ipin B3
*.opin adder_out3
*.opin Cout
*.ipin A0
x1 VDD VSS A0 adder_out0 B0 net1 VSS 1bit_adder
x2 VDD VSS A1 adder_out1 B1 net2 net1 1bit_adder
x3 VDD VSS A2 adder_out2 B2 net3 net2 1bit_adder
x4 VDD VSS A3 adder_out3 B3 Cout net3 1bit_adder
.ends


* expanding   symbol:  and/and2.sym # of pins=5
** sym_path: /home/halil/Desktop/design/xschem/and/and2.sym
** sch_path: /home/halil/Desktop/design/xschem/and/and2.sch
.subckt and2  VSS VDD A out B
*.ipin VDD
*.ipin A
*.ipin B
*.ipin VSS
*.opin out
XM1 net1 A net2 net2 sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 net1 A VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 net2 B VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 net1 B VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 out net1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 out net1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends


* expanding   symbol:  1bit_adder.sym # of pins=7
** sym_path: /home/halil/Desktop/design/xschem/1bit_adder.sym
** sch_path: /home/halil/Desktop/design/xschem/1bit_adder.sch
.subckt 1bit_adder  VDD VSS A adder_out B Cout Cin
*.ipin A
*.ipin B
*.iopin VDD
*.iopin VSS
*.ipin Cin
*.opin Cout
*.opin adder_out
x1 A B VDD VSS net1 xor2
x2 VSS VDD A net2 B and2
x3 VSS VDD net1 net3 Cin and2
x4 net1 Cin VDD VSS adder_out xor2
x5 net3 net2 VDD VSS Cout xor2
x6 net1 Cin VDD VSS adder_out xor2
.ends


* expanding   symbol:  xor2/xor2.sym # of pins=5
** sym_path: /home/halil/Desktop/design/xschem/xor2/xor2.sym
** sch_path: /home/halil/Desktop/design/xschem/xor2/xor2.sch
.subckt xor2  A B VDD VSS out
*.ipin A
*.ipin B
*.opin out
*.ipin VDD
*.ipin VSS
XM1 out notA net3 net3 sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 out B net1 net1 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 net3 notB VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 net1 notA VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 net4 A VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 out notB net4 net4 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM7 out A net2 net2 sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM8 net2 B VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM9 notA A VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM10 notA A VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM11 notB B VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM12 notB B VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
