** sch_path: /home/halil/Desktop/design/xschem/inv/inv_8bit.sch
**.subckt inv_8bit A0 A1 A2 A3 A4 A5 A6 A7 B0 B1 B2 B3 B4 B5 B6 B7 VDD VSS
*.ipin A0
*.ipin A1
*.ipin A2
*.ipin A3
*.ipin A4
*.ipin A5
*.ipin A6
*.ipin A7
*.opin B0
*.opin B1
*.opin B2
*.opin B3
*.opin B4
*.opin B5
*.opin B6
*.opin B7
*.ipin VDD
*.ipin VSS
x1 A0 VDD VSS B0 inverter
x2 A1 VDD VSS B1 inverter
x3 A2 VDD VSS B2 inverter
x4 A3 VDD VSS B3 inverter
x5 A4 VDD VSS B4 inverter
x6 A5 VDD VSS B5 inverter
x7 A6 VDD VSS B6 inverter
x8 A7 VDD VSS B7 inverter
**.ends

* expanding   symbol:  inv/inverter.sym # of pins=4
** sym_path: /home/halil/Desktop/design/xschem/inv/inverter.sym
** sch_path: /home/halil/Desktop/design/xschem/inv/inverter.sch
.subckt inverter  in Vdd Vss out
*.ipin in
*.iopin Vdd
*.iopin Vss
*.opin out
XM2 out in Vss Vss sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM11 out in Vdd Vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
