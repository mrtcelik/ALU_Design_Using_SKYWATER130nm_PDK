** sch_path: /home/halil/Desktop/design/xschem/or2_8bit.sch
**.subckt or2_8bit A0 Y0 B0 VDD VSS A1 B1 Y1 A2 B2 Y2 A3 B3 Y3 A4 B4 Y4 A5 B5 Y5 Y6 A6 B6 B7 A7 Y7
*.ipin A0
*.opin Y0
*.ipin B0
*.ipin VDD
*.ipin VSS
*.ipin A1
*.ipin B1
*.opin Y1
*.ipin A2
*.ipin B2
*.opin Y2
*.ipin A3
*.ipin B3
*.opin Y3
*.ipin A4
*.ipin B4
*.opin Y4
*.ipin A5
*.ipin B5
*.opin Y5
*.opin Y6
*.ipin A6
*.ipin B6
*.ipin B7
*.ipin A7
*.opin Y7
x1 VSS VDD A0 B0 Y0 or2
x2 VSS VDD A1 B1 Y1 or2
x3 VSS VDD A2 B2 Y2 or2
x4 VSS VDD A3 B3 Y3 or2
x5 VSS VDD A4 B4 Y4 or2
x6 VSS VDD A5 B5 Y5 or2
x7 VSS VDD A6 B6 Y6 or2
x8 VSS VDD A7 B7 Y7 or2
**.ends

* expanding   symbol:  or2.sym # of pins=5
** sym_path: /home/halil/Desktop/design/xschem/or2.sym
** sch_path: /home/halil/Desktop/design/xschem/or2.sch
.subckt or2  VSS VDD A B out
*.ipin A
*.ipin B
*.opin out
*.ipin VSS
*.ipin VDD
XM1 net2 B VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 net2 B net1 net1 sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 net1 A VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 net2 A VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 out net2 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 out net2 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
