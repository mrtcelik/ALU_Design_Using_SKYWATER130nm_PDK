** sch_path: /home/halil/Desktop/design/xschem/and2_8bit.sch
**.subckt and2_8bit A0 B0 VDD VSS Y0 A1 B1 Y1 A2 B2 Y2 A3 B3 Y3 A4 B4 Y4 A5 B5 Y5 A6 B6 Y6 A7 B7 Y7
*.ipin A0
*.ipin B0
*.ipin VDD
*.ipin VSS
*.opin Y0
*.ipin A1
*.ipin B1
*.opin Y1
*.ipin A2
*.ipin B2
*.opin Y2
*.ipin A3
*.ipin B3
*.opin Y3
*.ipin A4
*.ipin B4
*.opin Y4
*.ipin A5
*.ipin B5
*.opin Y5
*.ipin A6
*.ipin B6
*.opin Y6
*.ipin A7
*.ipin B7
*.opin Y7
x1 VSS VDD A0 Y0 B0 and2
x2 VSS VDD A1 Y1 B1 and2
x3 VSS VDD A2 Y2 B2 and2
x4 VSS VDD A3 Y3 B3 and2
x5 VSS VDD A4 Y4 B4 and2
x6 VSS VDD A5 Y5 B5 and2
x7 VSS VDD A6 Y6 B6 and2
x8 VSS VDD A7 Y7 B7 and2
**.ends

* expanding   symbol:  and2.sym # of pins=5
** sym_path: /home/halil/Desktop/design/xschem/and2.sym
** sch_path: /home/halil/Desktop/design/xschem/and2.sch
.subckt and2  VSS VDD A out B
*.ipin VDD
*.ipin A
*.ipin B
*.ipin VSS
*.opin out
XM1 net1 A net2 net2 sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 net1 A VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM3 net2 B VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM4 net1 B VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM5 out net1 VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM6 out net1 VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
