** sch_path: /home/halil/Desktop/design/xschem/hw4.sch
**.subckt hw4
XM2 clk3 Vdd net1 Vdd sky130_fd_pr__nfet_01v8 L=0.15 W=1.94 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM11 clk3 GND net1 GND sky130_fd_pr__pfet_01v8 L=0.15 W=4.76 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
R1 clk net1 750 m=1
V1 clk GND pulse(1.2 0 0 .1p .1p 50n 100n)
R2 net1 net2 750 m=1
R3 net2 clk2 750 m=1
R4 net2 clk1 750 m=1
C1 clk1 GND 200f m=1
C2 clk2 GND 200f m=1
C3 clk3 GND 200f m=1
C4 net2 GND 200f m=1
C5 net1 GND 200f m=1
V2 Vdd GND 1.2
**** begin user architecture code

** opencircuitdesign pdks install
.lib /usr/local/share/pdk/sky130B/libs.tech/ngspice/sky130.lib.spice tt_mm




.control
save all
tran 1n 200n
set color0=white

plot clk clk1+2 clk2+4 clk3+6
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
